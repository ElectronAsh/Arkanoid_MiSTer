
module source (
	source,
	probe);	

	output	[7:0]	source;
	input	[7:0]	probe;
endmodule
